 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity dp_ram_byte0 is
    port(clka : in std_logic;
    clkb : in std_logic;
    ena : in std_logic;
    enb : in std_logic;
    wea : in std_logic_vector(0 downto 0);
    web : in std_logic_vector(0 downto 0);
    addra : in std_logic_vector(8 downto 0);
    addrb : in std_logic_vector(8 downto 0);
    dia : in std_logic_vector(7 downto 0);
    dib : in std_logic_vector(7 downto 0);
    doa : out std_logic_vector(7 downto 0);
    dob : out std_logic_vector(7 downto 0));
end dp_ram_byte0;
architecture arch_dp_ram_byte0 of dp_ram_byte0 is
    type ram_type is array (511 downto 0) of std_logic_vector(7 downto 0);
    shared variable RAM : ram_type:= (
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"83",   
   X"06",   
   X"88",   
   X"09",   
   X"88",   
   X"06",   
   X"81",   
   X"fa",   
   X"6f",   
   X"e1",   
   X"4f",   
   X"b9",   
   X"1e",   
   X"7f",   
   X"da",   
   X"2f",   
   X"7f",   
   X"c8",   
   X"0a",   
   X"45",   
   X"79",   
   X"a4",   
   X"c8",   
   X"e3",   
   X"f6",   
   X"ff",   
   X"ff",   
   X"f6",   
   X"e2",   
   X"c4",   
   X"9b",   
   X"68",   
   X"29",   
   X"df",   
   X"89",   
   X"27",   
   X"ba",   
   X"3f",   
   X"b8",   
   X"24",   
   X"83",   
   X"d4",   
   X"18",   
   X"4f",   
   X"77",   
   X"91",   
   X"9d",   
   X"9a",   
   X"89",   
   X"6a",   
   X"3b",   
   X"fd",   
   X"b0",   
   X"54",   
   X"e9",   
   X"6e",   
   X"e4",   
   X"4a",   
   X"a1",   
   X"e8",   
   X"1f",   
   X"46",   
   X"5e",   
   X"66",   
   X"5e",   
   X"46",   
   X"1f",   
   X"e8",   
   X"a1",   
   X"4a",   
   X"e4",   
   X"6e",   
   X"e9",   
   X"54",   
   X"b0",   
   X"fd",   
   X"3b",   
   X"6a",   
   X"89",   
   X"9a",   
   X"9d",   
   X"91",   
   X"77",   
   X"4f",   
   X"18",   
   X"d4",   
   X"83",   
   X"24",   
   X"b8",   
   X"3f",   
   X"ba",   
   X"28",   
   X"89",   
   X"df",   
   X"29",   
   X"68",   
   X"9b",   
   X"c4",   
   X"e2",   
   X"f6",   
   X"ff",   
   X"ff",   
   X"f6",   
   X"e3",   
   X"c8",   
   X"a4",   
   X"79",   
   X"45",   
   X"0a",   
   X"c8",   
   X"7f",   
   X"2f",   
   X"da",   
   X"7f",   
   X"1f",   
   X"b9",   
   X"4f",   
   X"e1",   
   X"6f",   
   X"fa",   
   X"81",   
   X"06",   
   X"88",   
   X"09",   
   X"88",   
   X"06",   
   X"83",   
   X"00",   
   X"7c",   
   X"f9",   
   X"77",   
   X"f6",   
   X"77",   
   X"f9",   
   X"7e",   
   X"05",   
   X"90",   
   X"1e",   
   X"b0",   
   X"46",   
   X"e1",   
   X"80",   
   X"25",   
   X"d0",   
   X"80",   
   X"37",   
   X"f5",   
   X"ba",   
   X"87",   
   X"5b",   
   X"37",   
   X"1c",   
   X"09",   
   X"00",   
   X"00",   
   X"09",   
   X"1d",   
   X"3b",   
   X"64",   
   X"97",   
   X"d6",   
   X"20",   
   X"76",   
   X"d8",   
   X"46",   
   X"c0",   
   X"47",   
   X"db",   
   X"7c",   
   X"2b",   
   X"e7",   
   X"b1",   
   X"88",   
   X"6e",   
   X"62",   
   X"65",   
   X"76",   
   X"96",   
   X"c4",   
   X"02",   
   X"4f",   
   X"ab",   
   X"16",   
   X"91",   
   X"1b",   
   X"b5",   
   X"5e",   
   X"17",   
   X"e0",   
   X"b9",   
   X"a1",   
   X"99",   
   X"a1",   
   X"b9",   
   X"e0",   
   X"17",   
   X"5e",   
   X"b5",   
   X"1b",   
   X"91",   
   X"16",   
   X"ab",   
   X"4f",   
   X"02",   
   X"c4",   
   X"95",   
   X"76",   
   X"65",   
   X"62",   
   X"6e",   
   X"88",   
   X"b0",   
   X"e7",   
   X"2b",   
   X"7c",   
   X"db",   
   X"47",   
   X"c0",   
   X"45",   
   X"d7",   
   X"76",   
   X"20",   
   X"d6",   
   X"97",   
   X"64",   
   X"3b",   
   X"1d",   
   X"09",   
   X"ff",   
   X"ff",   
   X"09",   
   X"1b",   
   X"37",   
   X"5a",   
   X"86",   
   X"ba",   
   X"f5",   
   X"37",   
   X"80",   
   X"d0",   
   X"25",   
   X"80",   
   X"e0",   
   X"46",   
   X"b0",   
   X"1e",   
   X"90",   
   X"05",   
   X"7e",   
   X"f9",   
   X"76",   
   X"f6",   
   X"77",   
   X"f9",   
   X"7c"   
); 
 begin 
 process (CLKA) 
  begin 
  if (rising_edge(CLKA)) then 
   if ENA = '1' then 
    if WEA(0) = '1' then 
      RAM(conv_integer(ADDRA)) := DIA; 
    end if; 
   DOA <= RAM(conv_integer(ADDRA)); 
   end if; 
  end if; 
 end process; 
 process (CLKB) 
  begin 
   if (rising_edge(CLKB)) then 
    if ENB = '1' then 
      if WEB(0) = '1' then 
        RAM(conv_integer(ADDRB)) := DIB; 
      end if; 
    DOB <= RAM(conv_integer(ADDRB)); 
   end if; 
  end if; 
 end process; 
 end arch_dp_ram_byte0;  
