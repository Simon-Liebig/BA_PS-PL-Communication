 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity dp_ram_byte2 is
    port(clka : in std_logic;
    clkb : in std_logic;
    ena : in std_logic;
    enb : in std_logic;
    wea : in std_logic_vector(0 downto 0);
    web : in std_logic_vector(0 downto 0);
    addra : in std_logic_vector(8 downto 0);
    addrb : in std_logic_vector(8 downto 0);
    dia : in std_logic_vector(7 downto 0);
    dib : in std_logic_vector(7 downto 0);
    doa : out std_logic_vector(7 downto 0);
    dob : out std_logic_vector(7 downto 0));
end dp_ram_byte2;
architecture arch_dp_ram_byte2 of dp_ram_byte2 is
    type ram_type is array (511 downto 0) of std_logic_vector(7 downto 0);
    shared variable RAM : ram_type:= (
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"41",   
   X"c4",   
   X"47",   
   X"c9",   
   X"49",   
   X"c7",   
   X"44",   
   X"be",   
   X"35",   
   X"a9",   
   X"19",   
   X"85",   
   X"ec",   
   X"4f",   
   X"ad",   
   X"05",   
   X"58",   
   X"a4",   
   X"ea",   
   X"28",   
   X"60",   
   X"8f",   
   X"b7",   
   X"d7",   
   X"ee",   
   X"fc",   
   X"01",   
   X"fc",   
   X"ed",   
   X"d4",   
   X"b1",   
   X"83",   
   X"4a",   
   X"06",   
   X"b6",   
   X"5a",   
   X"f2",   
   X"7e",   
   X"fd",   
   X"70",   
   X"d5",   
   X"2d",   
   X"78",   
   X"b5",   
   X"e4",   
   X"06",   
   X"19",   
   X"1e",   
   X"14",   
   X"fb",   
   X"d4",   
   X"9e",   
   X"59",   
   X"04",   
   X"a1",   
   X"2d",   
   X"ab",   
   X"19",   
   X"77",   
   X"c6",   
   X"05",   
   X"35",   
   X"54",   
   X"64",   
   X"64",   
   X"54",   
   X"35",   
   X"05",   
   X"c6",   
   X"77",   
   X"19",   
   X"ab",   
   X"2e",   
   X"a1",   
   X"04",   
   X"59",   
   X"9e",   
   X"d4",   
   X"fb",   
   X"14",   
   X"1e",   
   X"19",   
   X"06",   
   X"e4",   
   X"b5",   
   X"78",   
   X"2d",   
   X"d5",   
   X"70",   
   X"fd",   
   X"7e",   
   X"f2",   
   X"5a",   
   X"b6",   
   X"06",   
   X"4a",   
   X"83",   
   X"b1",   
   X"d4",   
   X"ed",   
   X"fc",   
   X"01",   
   X"fc",   
   X"ee",   
   X"d7",   
   X"b7",   
   X"90",   
   X"60",   
   X"28",   
   X"ea",   
   X"a4",   
   X"58",   
   X"05",   
   X"ad",   
   X"4f",   
   X"ec",   
   X"85",   
   X"19",   
   X"a9",   
   X"35",   
   X"be",   
   X"44",   
   X"c8",   
   X"49",   
   X"c9",   
   X"47",   
   X"c4",   
   X"41",   
   X"be",   
   X"3b",   
   X"b8",   
   X"36",   
   X"b6",   
   X"38",   
   X"bb",   
   X"41",   
   X"ca",   
   X"57",   
   X"e6",   
   X"7a",   
   X"13",   
   X"b0",   
   X"52",   
   X"fa",   
   X"a7",   
   X"5b",   
   X"16",   
   X"d7",   
   X"9f",   
   X"70",   
   X"48",   
   X"28",   
   X"11",   
   X"03",   
   X"fe",   
   X"03",   
   X"12",   
   X"2b",   
   X"4e",   
   X"7c",   
   X"b5",   
   X"f9",   
   X"49",   
   X"a5",   
   X"0d",   
   X"81",   
   X"02",   
   X"8f",   
   X"2a",   
   X"d2",   
   X"87",   
   X"4a",   
   X"1b",   
   X"f9",   
   X"e6",   
   X"e2",   
   X"eb",   
   X"04",   
   X"2b",   
   X"61",   
   X"a6",   
   X"fb",   
   X"5e",   
   X"d2",   
   X"54",   
   X"e6",   
   X"88",   
   X"39",   
   X"fa",   
   X"ca",   
   X"ab",   
   X"9b",   
   X"9b",   
   X"ab",   
   X"ca",   
   X"fa",   
   X"39",   
   X"88",   
   X"e6",   
   X"54",   
   X"d1",   
   X"5e",   
   X"fb",   
   X"a6",   
   X"61",   
   X"2b",   
   X"04",   
   X"eb",   
   X"e1",   
   X"e6",   
   X"f9",   
   X"1b",   
   X"4a",   
   X"87",   
   X"d2",   
   X"2a",   
   X"8f",   
   X"02",   
   X"81",   
   X"0d",   
   X"a5",   
   X"49",   
   X"f9",   
   X"b5",   
   X"7c",   
   X"4e",   
   X"2b",   
   X"12",   
   X"03",   
   X"fe",   
   X"03",   
   X"11",   
   X"28",   
   X"48",   
   X"6f",   
   X"9f",   
   X"d7",   
   X"15",   
   X"5b",   
   X"a7",   
   X"fa",   
   X"52",   
   X"b0",   
   X"12",   
   X"7a",   
   X"e6",   
   X"56",   
   X"ca",   
   X"41",   
   X"bb",   
   X"37",   
   X"b6",   
   X"36",   
   X"b8",   
   X"3a",   
   X"be"   
); 
 begin 
 process (CLKA) 
  begin 
  if (rising_edge(CLKA)) then 
   if ENA = '1' then 
    if WEA(0) = '1' then 
      RAM(conv_integer(ADDRA)) := DIA; 
    end if; 
   DOA <= RAM(conv_integer(ADDRA)); 
   end if; 
  end if; 
 end process; 
 process (CLKB) 
  begin 
   if (rising_edge(CLKB)) then 
    if ENB = '1' then 
      if WEB(0) = '1' then 
        RAM(conv_integer(ADDRB)) := DIB; 
      end if; 
    DOB <= RAM(conv_integer(ADDRB)); 
   end if; 
  end if; 
 end process; 
 end arch_dp_ram_byte2;  
