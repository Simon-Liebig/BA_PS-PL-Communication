 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity dp_ram_byte3 is
    port(clka : in std_logic;
    clkb : in std_logic;
    ena : in std_logic;
    enb : in std_logic;
    wea : in std_logic_vector(0 downto 0);
    web : in std_logic_vector(0 downto 0);
    addra : in std_logic_vector(8 downto 0);
    addrb : in std_logic_vector(8 downto 0);
    dia : in std_logic_vector(7 downto 0);
    dib : in std_logic_vector(7 downto 0);
    doa : out std_logic_vector(7 downto 0);
    dob : out std_logic_vector(7 downto 0));
end dp_ram_byte3;
architecture arch_dp_ram_byte3 of dp_ram_byte3 is
    type ram_type is array (511 downto 0) of std_logic_vector(7 downto 0);
    shared variable RAM : ram_type:= (
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"00",   
   X"81",   
   X"83",   
   X"86",   
   X"88",   
   X"8b",   
   X"8d",   
   X"90",   
   X"92",   
   X"95",   
   X"97",   
   X"9a",   
   X"9c",   
   X"9e",   
   X"a1",   
   X"a3",   
   X"a6",   
   X"a8",   
   X"aa",   
   X"ac",   
   X"af",   
   X"b1",   
   X"b3",   
   X"b5",   
   X"b7",   
   X"b9",   
   X"bb",   
   X"be",   
   X"bf",   
   X"c1",   
   X"c3",   
   X"c5",   
   X"c7",   
   X"c9",   
   X"cb",   
   X"cc",   
   X"ce",   
   X"cf",   
   X"d1",   
   X"d2",   
   X"d4",   
   X"d5",   
   X"d7",   
   X"d8",   
   X"d9",   
   X"da",   
   X"dc",   
   X"dd",   
   X"de",   
   X"df",   
   X"df",   
   X"e0",   
   X"e1",   
   X"e2",   
   X"e3",   
   X"e3",   
   X"e4",   
   X"e4",   
   X"e5",   
   X"e5",   
   X"e5",   
   X"e6",   
   X"e6",   
   X"e6",   
   X"e6",   
   X"e6",   
   X"e6",   
   X"e6",   
   X"e6",   
   X"e5",   
   X"e5",   
   X"e5",   
   X"e4",   
   X"e4",   
   X"e3",   
   X"e3",   
   X"e2",   
   X"e1",   
   X"e0",   
   X"df",   
   X"df",   
   X"de",   
   X"dd",   
   X"dc",   
   X"da",   
   X"d9",   
   X"d8",   
   X"d7",   
   X"d5",   
   X"d4",   
   X"d2",   
   X"d1",   
   X"cf",   
   X"ce",   
   X"cc",   
   X"cb",   
   X"c9",   
   X"c7",   
   X"c5",   
   X"c3",   
   X"c1",   
   X"bf",   
   X"be",   
   X"bb",   
   X"b9",   
   X"b7",   
   X"b5",   
   X"b3",   
   X"b1",   
   X"af",   
   X"ac",   
   X"aa",   
   X"a8",   
   X"a6",   
   X"a3",   
   X"a1",   
   X"9e",   
   X"9c",   
   X"9a",   
   X"97",   
   X"95",   
   X"92",   
   X"90",   
   X"8d",   
   X"8b",   
   X"88",   
   X"86",   
   X"83",   
   X"81",   
   X"7e",   
   X"7c",   
   X"79",   
   X"77",   
   X"74",   
   X"72",   
   X"6f",   
   X"6d",   
   X"6a",   
   X"68",   
   X"65",   
   X"63",   
   X"61",   
   X"5e",   
   X"5c",   
   X"59",   
   X"57",   
   X"55",   
   X"53",   
   X"50",   
   X"4e",   
   X"4c",   
   X"4a",   
   X"48",   
   X"46",   
   X"44",   
   X"41",   
   X"40",   
   X"3e",   
   X"3c",   
   X"3a",   
   X"38",   
   X"36",   
   X"34",   
   X"33",   
   X"31",   
   X"30",   
   X"2e",   
   X"2d",   
   X"2b",   
   X"2a",   
   X"28",   
   X"27",   
   X"26",   
   X"25",   
   X"23",   
   X"22",   
   X"21",   
   X"20",   
   X"20",   
   X"1f",   
   X"1e",   
   X"1d",   
   X"1c",   
   X"1c",   
   X"1b",   
   X"1b",   
   X"1a",   
   X"1a",   
   X"1a",   
   X"19",   
   X"19",   
   X"19",   
   X"19",   
   X"19",   
   X"19",   
   X"19",   
   X"19",   
   X"1a",   
   X"1a",   
   X"1a",   
   X"1b",   
   X"1b",   
   X"1c",   
   X"1c",   
   X"1d",   
   X"1e",   
   X"1f",   
   X"20",   
   X"20",   
   X"21",   
   X"22",   
   X"23",   
   X"25",   
   X"26",   
   X"27",   
   X"28",   
   X"2a",   
   X"2b",   
   X"2d",   
   X"2e",   
   X"30",   
   X"31",   
   X"33",   
   X"34",   
   X"36",   
   X"38",   
   X"3a",   
   X"3c",   
   X"3e",   
   X"40",   
   X"41",   
   X"44",   
   X"46",   
   X"48",   
   X"4a",   
   X"4c",   
   X"4e",   
   X"50",   
   X"53",   
   X"55",   
   X"57",   
   X"59",   
   X"5c",   
   X"5e",   
   X"61",   
   X"63",   
   X"65",   
   X"68",   
   X"6a",   
   X"6d",   
   X"6f",   
   X"72",   
   X"74",   
   X"77",   
   X"79",   
   X"7c",   
   X"7e"   
); 
 begin 
 process (CLKA) 
  begin 
  if (rising_edge(CLKA)) then 
   if ENA = '1' then 
    if WEA(0) = '1' then 
      RAM(conv_integer(ADDRA)) := DIA; 
    end if; 
   DOA <= RAM(conv_integer(ADDRA)); 
   end if; 
  end if; 
 end process; 
 process (CLKB) 
  begin 
   if (rising_edge(CLKB)) then 
    if ENB = '1' then 
      if WEB(0) = '1' then 
        RAM(conv_integer(ADDRB)) := DIB; 
      end if; 
    DOB <= RAM(conv_integer(ADDRB)); 
   end if; 
  end if; 
 end process; 
 end arch_dp_ram_byte3;  
